//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Thu Dec 12 13:17:40 2024
// Version: v11.9 11.9.0.4
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// lzy_SD2
module lzy_SD2(
    // Inputs
    EI,
    I,
    // Outputs
    Y
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input        EI;
input  [7:0] I;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output [7:0] Y;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire         EI;
wire   [7:0] I;
wire   [0:0] lzy_74HC148_0_A0to0;
wire   [1:1] lzy_74HC148_0_A1to1;
wire   [2:2] lzy_74HC148_0_A2to2;
wire         lzy_74HC148_0_GS;
wire   [7:0] Y_net_0;
wire   [7:0] Y_net_1;
wire   [2:0] A_net_0;
wire   [3:0] A_net_1;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire         GND_net;
wire         VCC_net;
//--------------------------------------------------------------------
// Inverted Nets
//--------------------------------------------------------------------
wire         GS_OUT_PRE_INV0_0;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign GND_net    = 1'b0;
assign VCC_net    = 1'b1;
//--------------------------------------------------------------------
// Inversions
//--------------------------------------------------------------------
assign lzy_74HC148_0_GS = ~ GS_OUT_PRE_INV0_0;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign Y_net_1 = Y_net_0;
assign Y[7:0]  = Y_net_1;
//--------------------------------------------------------------------
// Slices assignments
//--------------------------------------------------------------------
assign lzy_74HC148_0_A0to0[0] = A_net_0[0:0];
assign lzy_74HC148_0_A1to1[1] = A_net_0[1:1];
assign lzy_74HC148_0_A2to2[2] = A_net_0[2:2];
//--------------------------------------------------------------------
// Concatenation assignments
//--------------------------------------------------------------------
assign A_net_1 = { 1'b0 , lzy_74HC148_0_A2to2[2] , lzy_74HC148_0_A1to1[1] , lzy_74HC148_0_A0to0[0] };
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------lzy_74HC148
lzy_74HC148 lzy_74HC148_0(
        // Inputs
        .EI ( EI ),
        .I  ( I ),
        // Outputs
        .GS ( GS_OUT_PRE_INV0_0 ),
        .EO (  ),
        .A  ( A_net_0 ) 
        );

//--------lzy_74HC4511
lzy_74HC4511 lzy_74HC4511_0(
        // Inputs
        .LE ( GND_net ),
        .BI ( lzy_74HC148_0_GS ),
        .LT ( VCC_net ),
        .A  ( A_net_1 ),
        // Outputs
        .Y  ( Y_net_0 ) 
        );


endmodule
