//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Sat Dec 28 10:01:08 2024
// Version: v11.9 11.9.0.4
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// lzy_SD1
module lzy_SD1(
    // Inputs
    A,
    B,
    C,
    // Outputs
    Y
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input  A;
input  B;
input  C;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output Y;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire         A;
wire         B;
wire         C;
wire         Y_net_0;
wire         Y_net_1;
wire   [1:0] S_net_0;
wire   [3:0] I_net_0;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire         GND_net;
//--------------------------------------------------------------------
// Inverted Nets
//--------------------------------------------------------------------
wire   [0:0] I_IN_POST_INV0_0;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign GND_net    = 1'b0;
//--------------------------------------------------------------------
// Inversions
//--------------------------------------------------------------------
assign I_IN_POST_INV0_0[0] = ~ A;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign Y_net_1 = Y_net_0;
assign Y       = Y_net_1;
//--------------------------------------------------------------------
// Concatenation assignments
//--------------------------------------------------------------------
assign S_net_0 = { B , C };
assign I_net_0 = { A , 1'b0 , 1'b0 , I_IN_POST_INV0_0[0] };
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------lzy_74HC153
lzy_74HC153 lzy_74HC153_0(
        // Inputs
        .E ( GND_net ),
        .S ( S_net_0 ),
        .I ( I_net_0 ),
        // Outputs
        .Y ( Y_net_0 ) 
        );


endmodule
