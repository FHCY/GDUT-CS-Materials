//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Mon Nov 13 18:26:07 2023
// Version: v11.9 11.9.0.4
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// cyq_SD2
module cyq_SD2(
    // Inputs
    EI,
    I,
    // Outputs
    Y
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input        EI;
input  [0:7] I;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output [6:0] Y;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire   [0:0] cyq_74HC148_0_A0to0;
wire   [1:1] cyq_74HC148_0_A1to1;
wire   [2:2] cyq_74HC148_0_A2to2;
wire         cyq_74HC148_0_GS;
wire         EI;
wire   [0:7] I;
wire   [6:0] Y_net_0;
wire   [6:0] Y_net_1;
wire   [2:0] A_net_0;
wire   [3:0] D_net_0;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire         GND_net;
wire         VCC_net;
//--------------------------------------------------------------------
// Inverted Nets
//--------------------------------------------------------------------
wire   [0:0] A_OUT_PRE_INV0_0;
wire   [1:1] A_OUT_PRE_INV1_0;
wire   [2:2] A_OUT_PRE_INV2_0;
wire         GS_OUT_PRE_INV3_0;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign GND_net    = 1'b0;
assign VCC_net    = 1'b1;
//--------------------------------------------------------------------
// Inversions
//--------------------------------------------------------------------
assign cyq_74HC148_0_A0to0[0] = ~ A_OUT_PRE_INV0_0[0];
assign cyq_74HC148_0_A1to1[1] = ~ A_OUT_PRE_INV1_0[1];
assign cyq_74HC148_0_A2to2[2] = ~ A_OUT_PRE_INV2_0[2];
assign cyq_74HC148_0_GS       = ~ GS_OUT_PRE_INV3_0;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign Y_net_1 = Y_net_0;
assign Y[6:0]  = Y_net_1;
//--------------------------------------------------------------------
// Slices assignments
//--------------------------------------------------------------------
assign A_OUT_PRE_INV0_0[0] = A_net_0[0:0];
assign A_OUT_PRE_INV1_0[1] = A_net_0[1:1];
assign A_OUT_PRE_INV2_0[2] = A_net_0[2:2];
//--------------------------------------------------------------------
// Concatenation assignments
//--------------------------------------------------------------------
assign D_net_0 = { 1'b0 , cyq_74HC148_0_A2to2[2] , cyq_74HC148_0_A1to1[1] , cyq_74HC148_0_A0to0[0] };
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------cyq_74HC148
cyq_74HC148 cyq_74HC148_0(
        // Inputs
        .EI ( EI ),
        .I  ( I ),
        // Outputs
        .A  ( A_net_0 ),
        .GS ( GS_OUT_PRE_INV3_0 ),
        .EO (  ) 
        );

//--------cyq_74HC4511
cyq_74HC4511 cyq_74HC4511_0(
        // Inputs
        .LE ( GND_net ),
        .BI ( cyq_74HC148_0_GS ),
        .LT ( VCC_net ),
        .D  ( D_net_0 ),
        // Outputs
        .Y  ( Y_net_0 ) 
        );


endmodule
