`timescale 1ns/1ns

module test_cyq_comb;

endmodule

