//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Mon Nov 20 15:26:12 2023
// Version: v11.9 11.9.0.4
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// cyq_SD1
module cyq_SD1(
    // Inputs
    A,
    B,
    C,
    // Outputs
    Y
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input  A;
input  B;
input  C;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output Y;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire         A;
wire         B;
wire         C;
wire         Y_net_0;
wire         Y_net_1;
wire   [1:0] S_net_0;
wire   [0:3] I_net_0;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire         GND_net;
//--------------------------------------------------------------------
// Inverted Nets
//--------------------------------------------------------------------
wire   [1:1] I_IN_POST_INV0_0;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign GND_net    = 1'b0;
//--------------------------------------------------------------------
// Inversions
//--------------------------------------------------------------------
assign I_IN_POST_INV0_0[1] = ~ A;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign Y_net_1 = Y_net_0;
assign Y       = Y_net_1;
//--------------------------------------------------------------------
// Concatenation assignments
//--------------------------------------------------------------------
assign S_net_0 = { B , C };
assign I_net_0 = { 1'b0 , I_IN_POST_INV0_0[1] , A , 1'b0 };
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------cyq_74HC153
cyq_74HC153 cyq_74HC153_0(
        // Inputs
        .S ( S_net_0 ),
        .I ( I_net_0 ),
        .E ( GND_net ),
        // Outputs
        .Y ( Y_net_0 ) 
        );


endmodule
