//////////////////////////////////////////////////////////////////////
// Created by SmartDesign Tue Dec 23 19:37:14 2025
// Version: v11.9 11.9.0.4
//////////////////////////////////////////////////////////////////////

`timescale 1ns / 100ps

// lly_SD1
module lly_SD1(
    // Inputs
    EI,
    I1,
    I2,
    // Outputs
    Y
);

//--------------------------------------------------------------------
// Input
//--------------------------------------------------------------------
input        EI;
input  [7:0] I1;
input  [7:0] I2;
//--------------------------------------------------------------------
// Output
//--------------------------------------------------------------------
output [7:0] Y;
//--------------------------------------------------------------------
// Nets
//--------------------------------------------------------------------
wire         AND2_1_Y;
wire         AND2_2_Y;
wire         AND2_3_Y;
wire         EI;
wire   [7:0] I1;
wire   [7:0] I2;
wire   [0:0] lly_74HC148_0_A0to0;
wire   [1:1] lly_74HC148_0_A1to1;
wire   [2:2] lly_74HC148_0_A2to2;
wire         lly_74HC148_0_EO;
wire         lly_74HC148_0_GS;
wire   [0:0] lly_74HC148_1_A0to0;
wire   [1:1] lly_74HC148_1_A1to1;
wire   [2:2] lly_74HC148_1_A2to2;
wire   [7:0] Y_net_0;
wire   [7:0] Y_net_1;
wire   [2:0] A_net_0;
wire   [2:0] A_net_1;
wire   [3:0] A_net_2;
//--------------------------------------------------------------------
// TiedOff Nets
//--------------------------------------------------------------------
wire         GND_net;
wire         VCC_net;
//--------------------------------------------------------------------
// Inverted Nets
//--------------------------------------------------------------------
wire         GS_OUT_PRE_INV0_0;
//--------------------------------------------------------------------
// Constant assignments
//--------------------------------------------------------------------
assign GND_net = 1'b0;
assign VCC_net = 1'b1;
//--------------------------------------------------------------------
// Inversions
//--------------------------------------------------------------------
assign lly_74HC148_0_GS = ~ GS_OUT_PRE_INV0_0;
//--------------------------------------------------------------------
// Top level output port assignments
//--------------------------------------------------------------------
assign Y_net_1 = Y_net_0;
assign Y[7:0]  = Y_net_1;
//--------------------------------------------------------------------
// Slices assignments
//--------------------------------------------------------------------
assign lly_74HC148_0_A0to0[0] = A_net_0[0:0];
assign lly_74HC148_0_A1to1[1] = A_net_0[1:1];
assign lly_74HC148_0_A2to2[2] = A_net_0[2:2];
assign lly_74HC148_1_A0to0[0] = A_net_1[0:0];
assign lly_74HC148_1_A1to1[1] = A_net_1[1:1];
assign lly_74HC148_1_A2to2[2] = A_net_1[2:2];
//--------------------------------------------------------------------
// Concatenation assignments
//--------------------------------------------------------------------
assign A_net_2 = { lly_74HC148_0_GS , AND2_3_Y , AND2_2_Y , AND2_1_Y };
//--------------------------------------------------------------------
// Component instances
//--------------------------------------------------------------------
//--------AND2
AND2 AND2_1(
        // Inputs
        .A ( lly_74HC148_0_A0to0 ),
        .B ( lly_74HC148_1_A0to0 ),
        // Outputs
        .Y ( AND2_1_Y ) 
        );

//--------AND2
AND2 AND2_2(
        // Inputs
        .A ( lly_74HC148_0_A1to1 ),
        .B ( lly_74HC148_1_A1to1 ),
        // Outputs
        .Y ( AND2_2_Y ) 
        );

//--------AND2
AND2 AND2_3(
        // Inputs
        .A ( lly_74HC148_0_A2to2 ),
        .B ( lly_74HC148_1_A2to2 ),
        // Outputs
        .Y ( AND2_3_Y ) 
        );

//--------lly_74HC148
lly_74HC148 lly_74HC148_0(
        // Inputs
        .EI ( EI ),
        .I  ( I1 ),
        // Outputs
        .A  ( A_net_0 ),
        .GS ( GS_OUT_PRE_INV0_0 ),
        .EO ( lly_74HC148_0_EO ) 
        );

//--------lly_74HC148
lly_74HC148 lly_74HC148_1(
        // Inputs
        .EI ( lly_74HC148_0_EO ),
        .I  ( I2 ),
        // Outputs
        .A  ( A_net_1 ),
        .GS (  ),
        .EO (  ) 
        );

//--------lly_74HC4511
lly_74HC4511 lly_74HC4511_0(
        // Inputs
        .LE ( GND_net ),
        .BI ( lly_74HC148_0_GS ),
        .LT ( VCC_net ),
        .A  ( A_net_2 ),
        // Outputs
        .Y  ( Y_net_0 ) 
        );


endmodule
